library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity sine_wave_generator is
    port (
        clk      : in STD_LOGIC;
        reset    : in STD_LOGIC;
        y :  IN  STD_LOGIC_VECTOR(9 DOWNTO 0);
		x :  IN  STD_LOGIC_VECTOR(9 DOWNTO 0);
        sine_out : out STD_LOGIC
    );
end sine_wave_generator;

architecture behavioral of sine_wave_generator is
    type sine_wave_array is array (0 to 599) of integer;
    constant sine_wave : sine_wave_array := (
        317, 322, 327, 332, 336, 341, 345, 349, 354, 357, 361, 365, 368, 372, 375, 378, 380, 383, 385, 388, 390, 392, 393, 395, 396, 397, 398, 399, 399, 400, 400, 400, 400, 399, 399, 398, 397, 396, 394, 393, 391, 389, 387, 384, 382, 379, 376, 373, 370, 367, 363, 359, 356, 352, 347, 343, 339, 334, 329, 325, 320, 315, 309, 304, 299, 293, 288, 282, 276, 271, 265, 259, 253, 247, 241, 234, 228, 222, 216, 210, 203, 197, 191, 185, 178, 172, 166, 160, 154, 148, 142, 136, 130, 124, 118, 113, 107, 102, 96, 91, 86, 81, 76, 71, 66, 62, 57, 53, 49, 45, 41, 37, 34, 30, 27, 24, 21, 18, 16, 13, 11, 9, 8, 6, 4, 3, 2, 1, 1, 0, 0, 0, 0, 0, 1, 2, 3, 4, 5, 7, 8, 10, 12, 14, 17, 19, 22, 25, 28, 31, 35, 39, 42, 46, 50, 55, 59, 63, 68, 73, 78, 83, 88, 93, 98, 104, 109, 115, 121, 126, 132, 138, 144, 150, 156, 162, 168, 175, 181, 187, 193, 200, 206, 212, 218, 225, 231, 237, 243, 249, 255, 261, 267, 273, 279, 284, 290, 296, 301, 306, 312, 317, 322, 327, 331, 336, 341, 345, 349, 353, 357, 361, 365, 368, 371, 375, 377, 380, 383, 385, 388, 390, 392, 393, 395, 396, 397, 398, 399, 399, 400, 400, 400, 400, 399, 399, 398, 397, 396, 394, 393, 391, 389, 387, 385, 382, 379, 376, 373, 370, 367, 363, 360, 356, 352, 348, 343, 339, 334, 330, 325, 320, 315, 310, 304, 299, 294, 288, 282, 277, 271, 265, 259, 253, 247, 241, 235, 229, 222, 216, 210, 204, 197, 191, 185, 179, 173, 166, 160, 154, 148, 142, 136, 130, 124, 119, 113, 107, 102, 96, 91, 86, 81, 76, 71, 66, 62, 57, 53, 49, 45, 41, 37, 34, 30, 27, 24, 21, 18, 16, 14, 11, 9, 8, 6, 5, 3, 2, 1, 1, 0, 0, 0, 0, 0, 1, 2, 3, 4, 5, 6, 8, 10, 12, 14, 17, 19, 22, 25, 28, 31, 35, 38, 42, 46, 50, 54, 59, 63, 68, 72, 77, 82, 87, 93, 98, 103, 109, 115, 120, 126, 132, 138, 144, 150, 156, 162, 168, 174, 181, 187, 193, 199, 205, 212, 218, 224, 230, 237, 243, 249, 255, 261, 267, 273, 278, 284, 290, 295, 301, 306, 311, 316, 321, 326, 331, 336, 340, 345, 349, 353, 357, 361, 364, 368, 371, 374, 377, 380, 383, 385, 387, 390, 391, 393, 395, 396, 397, 398, 399, 399, 400, 400, 400, 400, 399, 399, 398, 397, 396, 394, 393, 391, 389, 387, 385, 382, 380, 377, 374, 370, 367, 364, 360, 356, 352, 348, 344, 339, 335, 330, 325, 320, 315, 310, 305, 299, 294, 288, 283, 277, 271, 265, 259, 253, 247, 241, 235, 229, 223, 217, 210, 204, 198, 192, 185, 179, 173, 167, 161, 154, 148, 142, 136, 131, 125, 119, 113, 108, 102, 97, 92, 86, 81, 76, 71, 67, 62, 58, 53, 49, 45, 41, 38, 34, 31, 27, 24, 21, 19, 16, 14, 12, 10, 8, 6, 5, 3, 2, 1, 1, 0, 0, 0, 0, 0, 1, 2, 3, 4, 5, 6, 8, 10, 12, 14, 16, 19, 22, 25, 28, 31, 35, 38, 42, 46, 50, 54, 58, 63, 67, 72, 77, 82, 87, 92, 98, 103, 109, 114, 120, 126, 132, 137, 143, 149, 155, 162, 168, 174, 180, 186, 193, 199, 205, 211, 218, 224, 230, 236, 242, 248, 254, 260, 266, 272, 278, 284, 289, 295
    );
    signal sine_value : integer := 0;
    signal sine_out_tmp : std_logic := '0';
    signal x_int : integer := to_integer(signed(x));
    signal y_int : integer := to_integer(signed(y));
begin
    process(clk, reset, x_int, y_int)
    begin
        if reset = '1' then
            sine_out_tmp <= '0';
        elsif (clk'event and clk = '1') then
            if(x_int >= 0 and x_int <= 599) then
                sine_value <= sine_wave(x_int);
                -- verifica se ta em cima da senoide
                if (y_int = sine_value) then
                    sine_out_tmp <= '1';
                else
                    sine_out_tmp <= '0';
                end if;
            else
                sine_out_tmp <= '0';
            end if;
        end if;
    end process;

    sine_out <= sine_out_tmp;
end behavioral;

-- Copyright (C) 2018  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.

-- Generated by Quartus Prime Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition
-- Created on Tue Apr 16 18:33:21 2024

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY robo_linha IS
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        sensorD : IN STD_LOGIC := '0';
        sensorE : IN STD_LOGIC := '0';
        timeout : IN STD_LOGIC := '0';
        velMotorD : OUT STD_LOGIC;
        velMotorE : OUT STD_LOGIC;
        esquerda : OUT STD_LOGIC;
        direita : OUT STD_LOGIC;
        perdido : OUT STD_LOGIC
    );
END robo_linha;

ARCHITECTURE BEHAVIOR OF robo_linha IS
    TYPE type_fstate IS (reto,virandoDireita,virandoEsquerda,parado,perdeuDireita,perdeuEsquerda);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,sensorD,sensorE,timeout)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= parado;
            velMotorD <= '0';
            velMotorE <= '0';
            esquerda <= '0';
            direita <= '0';
            perdido <= '0';
        ELSE
            velMotorD <= '0';
            velMotorE <= '0';
            esquerda <= '0';
            direita <= '0';
            perdido <= '0';
            CASE fstate IS
                WHEN reto =>
                    IF ((NOT((sensorE = '1')) AND (sensorD = '1'))) THEN
                        reg_fstate <= virandoDireita;
                    ELSIF (((sensorE = '1') AND NOT((sensorD = '1')))) THEN
                        reg_fstate <= virandoEsquerda;
                    ELSIF ((NOT((sensorE = '1')) AND NOT((sensorD = '1')))) THEN
                        reg_fstate <= parado;
                    ELSE
                        reg_fstate <= reto;
                    END IF;

                    esquerda <= '1';

                    velMotorE <= '1';

                    velMotorD <= '1';

                    perdido <= '0';

                    direita <= '1';
                WHEN virandoDireita =>
                    IF (((sensorE = '1') AND (sensorD = '1'))) THEN
                        reg_fstate <= reto;
                    ELSIF ((NOT((sensorE = '1')) AND NOT((sensorD = '1')))) THEN
                        reg_fstate <= perdeuDireita;
                    ELSE
                        reg_fstate <= virandoDireita;
                    END IF;

                    esquerda <= '0';

                    velMotorE <= '1';

                    velMotorD <= '0';

                    perdido <= '0';

                    direita <= '1';
                WHEN virandoEsquerda =>
                    IF (((sensorE = '1') AND (sensorD = '1'))) THEN
                        reg_fstate <= reto;
                    ELSIF ((NOT((sensorE = '1')) AND NOT((sensorD = '1')))) THEN
                        reg_fstate <= perdeuEsquerda;
                    ELSE
                        reg_fstate <= virandoEsquerda;
                    END IF;

                    esquerda <= '1';

                    velMotorE <= '0';

                    velMotorD <= '1';

                    perdido <= '0';

                    direita <= '0';
                WHEN parado =>
                    IF (((sensorE = '1') AND (sensorD = '1'))) THEN
                        reg_fstate <= reto;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= parado;
                    END IF;

                    esquerda <= '0';

                    velMotorE <= '0';

                    velMotorD <= '0';

                    perdido <= '0';

                    direita <= '0';
                WHEN perdeuDireita =>
                    IF ((((sensorE = '1') AND NOT((sensorD = '1'))) AND NOT((timeout = '1')))) THEN
                        reg_fstate <= virandoEsquerda;
                    ELSIF (((NOT((sensorE = '1')) AND NOT((sensorD = '1'))) AND NOT((timeout = '1')))) THEN
                        reg_fstate <= perdeuDireita;
                    ELSIF ((timeout = '1')) THEN
                        reg_fstate <= parado;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= perdeuDireita;
                    END IF;

                    velMotorE <= '0';

                    velMotorD <= '1';

                    perdido <= '1';
                WHEN perdeuEsquerda =>
                    IF (((NOT((sensorE = '1')) AND (sensorD = '1')) AND NOT((timeout = '1')))) THEN
                        reg_fstate <= virandoDireita;
                    ELSIF (((NOT((sensorE = '1')) AND NOT((sensorD = '1'))) AND NOT((timeout = '1')))) THEN
                        reg_fstate <= perdeuEsquerda;
                    ELSIF ((timeout = '1')) THEN
                        reg_fstate <= parado;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= perdeuEsquerda;
                    END IF;

                    velMotorE <= '1';

                    velMotorD <= '0';

                    perdido <= '1';
                WHEN OTHERS => 
                    velMotorD <= 'X';
                    velMotorE <= 'X';
                    esquerda <= 'X';
                    direita <= 'X';
                    perdido <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;

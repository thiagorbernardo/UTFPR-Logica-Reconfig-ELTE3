-- Copyright (C) 2018  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.


-- Generated by Quartus Prime Version 18.1 (Build Build 625 09/12/2018)
-- Created on Tue Apr 16 16:52:35 2024

robo_linha robo_linha_inst
(
	.clock(clock_sig) ,	// input  clock_sig
	.reset(reset_sig) ,	// input  reset_sig
	.sensorD(sensorD_sig) ,	// input  sensorD_sig
	.sensorE(sensorE_sig) ,	// input  sensorE_sig
	.timeout(timeout_sig) ,	// input  timeout_sig
	.velMotorD(velMotorD_sig) ,	// output  velMotorD_sig
	.velMotorE(velMotorE_sig) ,	// output  velMotorE_sig
	.esquerda(esquerda_sig) ,	// output  esquerda_sig
	.direita(direita_sig) ,	// output  direita_sig
	.perdido(perdido_sig) 	// output  perdido_sig
);


counter_inst : counter PORT MAP (
		clock	 => clock_sig,
		q	 => q_sig
	);

-- Copyright (C) 2018  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.

-- Generated by Quartus Prime Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition
-- Created on Tue Apr 25 12:09:24 2023

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY atividade1 IS
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        sensordir : IN STD_LOGIC := '0';
        sensoresq : IN STD_LOGIC := '0';
        velmotoresq : OUT STD_LOGIC;
        velmotordir : OUT STD_LOGIC;
        state1 : OUT STD_LOGIC;
        state0 : OUT STD_LOGIC
    );
END atividade1;

ARCHITECTURE BEHAVIOR OF atividade1 IS
    TYPE type_fstate IS (parado,esquerda,direita,reto);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,sensordir,sensoresq)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= parado;
            velmotoresq <= '0';
            velmotordir <= '0';
            state1 <= '0';
            state0 <= '0';
        ELSE
            velmotoresq <= '0';
            velmotordir <= '0';
            state1 <= '0';
            state0 <= '0';
            CASE fstate IS
                WHEN parado =>
                    IF (((sensoresq = '1') AND (sensordir = '1'))) THEN
                        reg_fstate <= reto;
                    ELSE
                        reg_fstate <= parado;
                    END IF;

                    state0 <= '0';

                    state1 <= '0';

                    velmotordir <= '0';

                    velmotoresq <= '0';
                WHEN esquerda =>
                    IF (((sensoresq = '1') AND (sensordir = '1'))) THEN
                        reg_fstate <= reto;
                    ELSIF ((NOT((sensoresq = '1')) AND NOT((sensordir = '1')))) THEN
                        reg_fstate <= parado;
                    ELSE
                        reg_fstate <= esquerda;
                    END IF;

                    state0 <= '1';

                    state1 <= '0';

                    velmotordir <= '1';

                    velmotoresq <= '0';
                WHEN direita =>
                    IF (((sensoresq = '1') AND (sensordir = '1'))) THEN
                        reg_fstate <= reto;
                    ELSIF ((NOT((sensoresq = '1')) AND NOT((sensordir = '1')))) THEN
                        reg_fstate <= parado;
                    ELSE
                        reg_fstate <= direita;
                    END IF;

                    state0 <= '0';

                    state1 <= '1';

                    velmotordir <= '0';

                    velmotoresq <= '1';
                WHEN reto =>
                    IF ((NOT((sensoresq = '1')) AND NOT((sensordir = '1')))) THEN
                        reg_fstate <= parado;
                    ELSIF ((NOT((sensoresq = '1')) AND (sensordir = '1'))) THEN
                        reg_fstate <= direita;
                    ELSIF (((sensoresq = '1') AND NOT((sensordir = '1')))) THEN
                        reg_fstate <= esquerda;
                    ELSE
                        reg_fstate <= reto;
                    END IF;

                    state0 <= '1';

                    state1 <= '1';

                    velmotordir <= '1';

                    velmotoresq <= '1';
                WHEN OTHERS => 
                    velmotoresq <= 'X';
                    velmotordir <= 'X';
                    state1 <= 'X';
                    state0 <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
